library IEEE;
use IEEE.STD_LOGIC_1164.all;
-- Entidade sem portos
entity DrinksFSM_Tb is
end DrinksFSM_Tb;


architecture Stimulus of DrinksFSM_Tb is
 -- Sinais para ligar às entradas da UUT
signal s_reset : std_logic;
signal s_clk : std_logic;
signal s_coin_20 : std_logic;
signal s_coin_50 : std_logic;

 -- Sinal para ligar às saídas da UUT
signal s_drinks : std_logic;



begin
 -- Instanciação da Unit Under Test (UUT)
 uut: entity work.DrinksFSM(Behavioral)
 port map(reset => s_reset,
			 clk => s_clk,
			coin_20 => s_coin_20,
			coin_50 => s_coin_20,
			drinks => s_drinks);
		
	
------- process clock
clock_proc : process

begin
s_clk <= '0'; wait for 50 ns;
s_clk <='1'; wait for 50 ns;
end process;
 --Process stim
 
 stim_proc : process

 begin

 s_reset <= '1';
 s_coin_20 <= '0';
 s_coin_50 <= '0';
 
wait for 325 ns;
s_reset <= '0';

wait for 30 ns;
s_coin_20 <='1';
s_coin_50 <= '0';
 
 wait for 600 ns;
 
 s_reset<= '1';
 
 wait for 110 ns;
 s_reset <= '0';
 s_coin_20 <= '0';
 s_coin_50 <= '1';
 wait for 200 ns;
s_reset <= '1';


 wait for 100 ns;
 s_reset <= '0';
 s_coin_20 <= '1';
 s_coin_50 <= '0';
 
  wait for 100 ns;
 s_reset <= '0';
 s_coin_20 <= '0';
 s_coin_50 <= '0';
 
 
 wait for 125 ns;
 s_coin_20 <='0';
 s_coin_50<='0';

 end process;
end Stimulus; 