use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

